// ------------------------------------------------------------------------- 
// File name    : AHB_UVC_defines.sv
// Title        : AHB_UVC defines
// Project      : AHB_UVC
// Created On   : 2024-02-07
// Developers   : 
// -------------------------------------------------------------------------

`define ADDR_WIDTH 8

