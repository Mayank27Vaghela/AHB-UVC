`ifndef AHB_UVC_PKG_SV
`define AHB_UVC_PKG_SV
package AHB_UVC_package;
   
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import AHB_UVC_master_package::*;
  import AHB_UVC_slave_package::*;
  import AHB_UVC_env_package::*;
  import AHB_UVC_test_package::*;

endpackage : AHB_UVC_package
`endif /** AHB_UVC_PKG*/
